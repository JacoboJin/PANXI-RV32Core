`timescale 1ns/1ps


`define DATA_WIDTH  = 32